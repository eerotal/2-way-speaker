Two-way speaker crossover filter

* Visaton W-170S model
.subckt W170S 1 2
RS 1 2 5.9
LS 2 3 1.2m
.ends

* Visaton SC-10N model
.subckt SC10N 1 2
RS 1 2 6.9
LS 2 3 0.04m
.ends


* Low-pass filter section
V1 GND in dc 0 ac { 14*1.414 }
L1 in L1_2 1m
C2 L1_2 GND 6.8u
R1 L1_2 R1_2 8.2
L3 L1_2 R1_2 1m
R4 R1_2 R4_2 8.2
VS_R4 R4_2 VS_R4_2 0
C4 VS_R4_2 GND 22u
XWOOFER R1_2 WOOFER_OUT W170S
VS_WOOFER WOOFER_OUT GND 0

* High-pass filter
C1 in C1_2 6.8u
L2 C1_2 GND 0.47m
C3 C1_2 C3_2 10u
R3 C3_2 R3_2 4.1
VS_R3 R3_2 VS_R3_2 0
R5 VS_R3_2 R5_2 4.1
VS_R5 R5_2 GND 0
XTWEETER VS_R3_2 TWEETER_OUT SC10N
VS_TWEETER TWEETER_OUT GND 0

* Simulation parameters.
.control
ac dec 100 15 10k

* Setup plot export options.
set hcopydevtype = postscript
set hcopypscolor = 1

* Plot resistor powers.
let R1_pwr = (v(L1_2) - v(R1_2))*i(VS_WOOFER)
let R4_pwr = (v(R4_2) - v(R1_2))*i(VS_R4)
let R3_pwr = (v(C3_2) - v(R3_2))*i(VS_R3)
let R5_pwr = (v(VS_R3_2) - v(R5_2))*i(VS_R5)
hardcopy r_pwr.ps R1_pwr R4_pwr R3_pwr R5_pwr ylabel 'Power (W)' xlabel 'Frequency' title 'Resistor power dissipation'

* Plot speaker powers.
let tweeter_pwr = (v(VS_R3_2) - v(TWEETER_OUT))*i(VS_TWEETER)
let woofer_pwr = (v(R1_2) - v(WOOFER_OUT))*i(VS_WOOFER)
hardcopy spk_pwr.ps tweeter_pwr woofer_pwr ylabel 'Power (W)' xlabel 'Frequency' title 'Driver power dissipation'

* Plot input power.
let input_pwr = v(in)*i(V1)
hardcopy in_pwr.ps input_pwr ylabel 'Power (W)' xlabel 'Frequency' title 'Input power'

* Plot voltage gains at speaker inputs.
let Vg_woofer = v(R1_2)/v(in)
let Vg_tweeter = v(R3_2)/v(in)
hardcopy gain.ps vdb(Vg_woofer) vdb(Vg_tweeter) ylabel 'Voltage gain (dB)' xlabel 'Frequency' title 'Voltage gain at speaker inputs'
.endc

.end

